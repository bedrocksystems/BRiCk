(*
 * Copyright (C) BedRock Systems Inc. 2019 Gregory Malecha
 *
 * SPDX-License-Identifier:AGPL-3.0-or-later
 *)

(** this module provides a denotational/axiomatic semantics to c++ compilation
    units.
 *)
From Coq.Classes Require Import
     RelationClasses Morphisms DecidableClass.

Require Import Coq.Lists.List.
Require Import Coq.Lists.List.
Require Import Coq.Strings.String.
Require Import Coq.ZArith.BinInt.
Require Import Coq.micromega.Lia.

From bedrock Require Import IrisBridge.
Require Import bedrock.lang.cpp.ast.
From bedrock.lang.cpp Require Import
     semantics logic.pred logic.path_pred logic.heap_pred.
From bedrock.lang.cpp Require Import logic.wp.
Require Import iris.proofmode.tactics.

Import ChargeNotation.

Section with_cpp.
  Context `{Σ : cpp_logic ti} {resolve:genv}.

  Set Default Proof Using "Σ resolve".

  Local Notation _global := (@_global resolve) (only parsing).
  Local Notation code_at := (@code_at _ Σ resolve) (only parsing).
  Local Notation method_at := (@method_at _ Σ resolve) (only parsing).
  Local Notation ctor_at := (@ctor_at _ Σ resolve) (only parsing).
  Local Notation dtor_at := (@dtor_at _ Σ resolve) (only parsing).
  Local Notation _field := (@_field resolve) (only parsing).
  Local Notation _super := (@_super resolve) (only parsing).
  Local Notation _sub := (@_sub resolve) (only parsing).

  Definition denoteSymbol (n : obj_name) (o : ObjValue) : mpred :=
    Exists a, _global n &~ a **
    match o with
    | Ovar _ e => empSP
    | Ofunction f =>
      match f.(f_body) return mpred with
      | None => empSP
      | Some body => code_at f a
      end
    | Omethod m =>
      match m.(m_body) return mpred with
      | None => emp
      | Some body =>
        method_at m a
      end
    | Oconstructor c =>
      match c.(c_body) return mpred with
      | None => empSP
      | Some body => ctor_at c a
      end
    | Odestructor d =>
      match d.(d_body) return mpred with
      | None => empSP
      | Some body => dtor_at d a
      end
    end.

  Global Instance: Persistent (denoteSymbol n o).
  Proof using .
    rewrite /denoteSymbol; destruct o; simpl; red.
    - iIntros "#H"; iModIntro; iFrame "#".
    - iIntros "#H"; iModIntro; iFrame "#".
    - iIntros "#H"; iModIntro; iFrame "#".
    - iIntros "#H"; iModIntro; iFrame "#".
    - iIntros "#H"; iModIntro; iFrame "#".
  Qed.

  Global Instance: Affine (denoteSymbol n o).
  Proof using . refine _. Qed.

  Definition initSymbol (n : obj_name) (o : ObjValue) : mpred :=
    Exists a, _global n &~ a **
    match o with
    | Ovar t (Some e) =>
      ltrue (*
      Exists Q : FreeTemps -> mpred,
      □ (_at (_eq a) (uninitR (resolve:=resolve) t 1) -*
         Forall ρ ti, wp_init (resolve:=resolve) ti ρ t (Vptr a) e Q) ** Q empSP
*)
      (* ^^ todo(gmm): static initialization is not yet supported *)
    | Ovar t None =>
      _at (_eq a) (uninitR (resolve:=resolve) t 1)
    | _ => empSP
    end.

  Definition denoteModule_def (d : compilation_unit) : mpred :=
    ([∗map] on ↦ o ∈ d.(symbols), denoteSymbol on o)%I **
    [| module_le d resolve.(genv_cu) |].
  Definition denoteModule_aux : seal (@denoteModule_def). by eexists. Qed.
  Definition denoteModule := denoteModule_aux.(unseal).
  Definition denoteModule_eq : @denoteModule = _ := denoteModule_aux.(seal_eq).

  Global Instance: Persistent (denoteModule module).
  Proof.
    red. rewrite denoteModule_eq /denoteModule_def; intros.
    iIntros "[#M #H]"; iFrame "#".
  Qed.

  Global Instance: Affine (denoteModule module).
  Proof using . refine _. Qed.

End with_cpp.

Arguments denoteModule _ : simpl never.
